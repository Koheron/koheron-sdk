`timescale 1 ns / 1 ps

module pdm_tb();
  parameter NBITS = 10;
 
  reg                       clk;
  reg                       rst;
  reg [NBITS-1:0]           data_in;
  wire                      pdm_out;
  wire [NBITS-1:0]          pdm_error;

  pdm # (
    .NBITS(NBITS)
  )
  DUT (
    .clk(clk),
    .rst(rst),
    .data_in(data_in),
    .pdm_out(pdm_out),
    .pdm_error(pdm_error)
  );

  parameter CLK_PERIOD = 8;

  initial begin
    clk = 1;
    rst = 1;
    data_in = 120;
    #(10*CLK_PERIOD)
    rst = 0;
    #(1000*CLK_PERIOD)
    data_in = 500;
    #(1000*CLK_PERIOD)
    data_in = 900;    
    #(100000*CLK_PERIOD)
    $finish;
  end

  always #(CLK_PERIOD/2) clk = ~clk;

endmodule
